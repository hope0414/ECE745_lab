14 uid=262235
20 atime=1548446481
